module day_12_solver (
    m_tready,
    s_tdata,
    clear,
    clock,
    s_tvalid,
    s_tready,
    m_tvalid,
    m_tlast,
    m_tdata
);

    input m_tready;
    input [7:0] s_tdata;
    input clear;
    input clock;
    input s_tvalid;
    output s_tready;
    output m_tvalid;
    output m_tlast;
    output [7:0] m_tdata;

    wire _99;
    wire _194;
    wire _195;
    wire _196;
    wire _197;
    wire _102;
    wire _103;
    reg _199;
    wire _1;
    reg _100;
    wire _204;
    wire _205;
    wire _206;
    wire _207;
    wire _202;
    wire _203;
    reg _208;
    wire _2;
    reg _201;
    wire _210;
    wire [6:0] _209;
    wire [7:0] _211;
    wire _213;
    wire _214;
    wire _1367;
    wire [3:0] _84;
    wire _7;
    wire [3:0] _1364;
    wire [3:0] _1363;
    wire [3:0] _1359;
    wire [3:0] _1360;
    wire [3:0] _1361;
    wire [3:0] _1362;
    wire [3:0] _212;
    wire [3:0] _1357;
    wire [3:0] _1358;
    wire [3:0] _198;
    wire [3:0] _104;
    wire _1353;
    wire _1354;
    wire [15:0] _1349;
    wire [15:0] _1345;
    wire [7:0] _1340;
    wire [7:0] _1339;
    wire [15:0] _1341;
    wire [11:0] _1335;
    wire [15:0] _1337;
    wire [1:0] _1332;
    wire [13:0] _1331;
    wire [15:0] _1333;
    wire [15:0] _1329;
    wire _1327;
    wire [15:0] _1330;
    wire _1326;
    wire [15:0] _1334;
    wire _1325;
    wire [15:0] _1338;
    wire _1324;
    wire [15:0] _1342;
    wire [4:0] _1322;
    wire _1323;
    wire [15:0] _1344;
    wire [15:0] _1346;
    wire [15:0] _1347;
    wire [15:0] _1348;
    wire _1350;
    wire _1351;
    wire _242;
    wire gnd;
    wire _240;
    wire vdd;
    reg _243;
    wire _8;
    wire [15:0] _629;
    wire [15:0] _630;
    wire _241;
    wire [15:0] _631;
    wire [7:0] _623;
    wire [15:0] _625;
    wire [11:0] _619;
    wire [15:0] _621;
    wire [13:0] _615;
    wire [15:0] _617;
    wire [14:0] _611;
    wire [15:0] _613;
    wire [3:0] _604;
    wire [3:0] _602;
    reg [3:0] _606;
    wire [3:0] _598;
    wire [3:0] _597;
    reg [3:0] _601;
    reg [3:0] _596;
    reg [3:0] _591;
    reg [3:0] _586;
    reg [3:0] _581;
    reg [3:0] _576;
    reg [3:0] _571;
    reg [3:0] _607;
    reg [3:0] _565;
    reg [3:0] _560;
    reg [3:0] _555;
    reg [3:0] _550;
    reg [3:0] _545;
    reg [3:0] _540;
    reg [3:0] _535;
    wire [3:0] _527;
    reg [3:0] _530;
    reg [3:0] _566;
    wire [3:0] _521;
    reg [3:0] _524;
    wire [3:0] _516;
    reg [3:0] _519;
    reg [3:0] _514;
    reg [3:0] _509;
    reg [3:0] _504;
    reg [3:0] _499;
    reg [3:0] _494;
    reg [3:0] _489;
    reg [3:0] _525;
    reg [3:0] _483;
    reg [3:0] _478;
    reg [3:0] _473;
    reg [3:0] _468;
    reg [3:0] _463;
    reg [3:0] _458;
    reg [3:0] _453;
    reg [3:0] _448;
    reg [3:0] _484;
    reg [3:0] _442;
    wire [3:0] _436;
    reg [3:0] _437;
    reg [3:0] _432;
    reg [3:0] _427;
    reg [3:0] _422;
    reg [3:0] _417;
    reg [3:0] _412;
    reg [3:0] _407;
    reg [3:0] _443;
    reg [3:0] _401;
    reg [3:0] _396;
    reg [3:0] _391;
    reg [3:0] _386;
    reg [3:0] _381;
    reg [3:0] _376;
    reg [3:0] _371;
    wire [1:0] _361;
    reg [3:0] _366;
    reg [2:0] _359;
    wire [2:0] _360;
    reg [3:0] _402;
    reg [2:0] _357;
    wire [2:0] _265;
    reg [2:0] _268;
    wire [2:0] _269;
    reg [2:0] _271;
    wire [2:0] _9;
    reg [2:0] _266;
    reg [2:0] _275;
    wire [2:0] _276;
    reg [2:0] _277;
    wire [2:0] _10;
    reg [2:0] _273;
    reg [2:0] _281;
    wire [2:0] _282;
    reg [2:0] _283;
    wire [2:0] _11;
    reg [2:0] _279;
    reg [2:0] _287;
    wire [2:0] _288;
    reg [2:0] _289;
    wire [2:0] _12;
    reg [2:0] _285;
    reg [2:0] _293;
    wire [2:0] _294;
    reg [2:0] _295;
    wire [2:0] _13;
    reg [2:0] _291;
    reg [2:0] _299;
    wire [2:0] _300;
    reg [2:0] _301;
    wire [2:0] _14;
    reg [2:0] _297;
    reg [2:0] _305;
    wire [2:0] _306;
    reg [2:0] _307;
    wire [2:0] _15;
    reg [2:0] _303;
    reg [2:0] _311;
    wire [2:0] _312;
    reg [2:0] _313;
    wire [2:0] _16;
    reg [2:0] _309;
    reg [2:0] _317;
    wire [2:0] _318;
    reg [2:0] _319;
    wire [2:0] _17;
    reg [2:0] _315;
    reg [2:0] _323;
    wire [2:0] _324;
    reg [2:0] _325;
    wire [2:0] _18;
    reg [2:0] _321;
    reg [2:0] _329;
    wire [2:0] _330;
    reg [2:0] _331;
    wire [2:0] _19;
    reg [2:0] _327;
    reg [2:0] _335;
    wire [2:0] _336;
    reg [2:0] _337;
    wire [2:0] _20;
    reg [2:0] _333;
    reg [2:0] _356;
    wire [2:0] _358;
    reg [3:0] _608;
    wire [11:0] _355;
    wire [15:0] _609;
    wire _352;
    wire [2:0] _350;
    wire _351;
    wire _353;
    wire [15:0] _610;
    wire _349;
    wire [15:0] _614;
    wire _348;
    wire [15:0] _618;
    wire _347;
    wire [15:0] _622;
    reg [7:0] _343;
    wire [7:0] _344;
    wire [3:0] _345;
    wire _346;
    wire [15:0] _626;
    wire [15:0] _627;
    wire _239;
    wire [15:0] _628;
    reg [15:0] _632;
    wire [15:0] _21;
    reg [15:0] _340[0:15];
    wire _232;
    wire _230;
    wire _229;
    wire _231;
    wire _233;
    wire [2:0] _236;
    wire [4:0] _228;
    wire [7:0] _237;
    reg [7:0] _226;
    wire [7:0] _640;
    wire [7:0] _641;
    reg [7:0] _643;
    wire [7:0] _644;
    wire [7:0] _645;
    wire [7:0] _646;
    reg [7:0] _637;
    wire [7:0] _638;
    wire [7:0] _639;
    reg [7:0] _647;
    wire [7:0] _22;
    reg [7:0] _185;
    wire [7:0] _654;
    reg [7:0] _656;
    wire [7:0] _657;
    wire [7:0] _658;
    wire [7:0] _659;
    reg [7:0] _650;
    wire [7:0] _651;
    wire [7:0] _652;
    reg [7:0] _660;
    wire [7:0] _23;
    reg [7:0] _183;
    wire [7:0] _667;
    reg [7:0] _669;
    wire [7:0] _670;
    wire [7:0] _671;
    wire [7:0] _672;
    reg [7:0] _663;
    wire [7:0] _664;
    wire [7:0] _665;
    reg [7:0] _673;
    wire [7:0] _24;
    reg [7:0] _181;
    wire [7:0] _680;
    reg [7:0] _682;
    wire [7:0] _683;
    wire [7:0] _684;
    wire [7:0] _685;
    reg [7:0] _676;
    wire [7:0] _677;
    wire [7:0] _678;
    reg [7:0] _686;
    wire [7:0] _25;
    reg [7:0] _179;
    wire [7:0] _693;
    reg [7:0] _695;
    wire [7:0] _696;
    wire [7:0] _697;
    wire [7:0] _698;
    reg [7:0] _689;
    wire [7:0] _690;
    wire [7:0] _691;
    reg [7:0] _699;
    wire [7:0] _26;
    reg [7:0] _177;
    wire [7:0] _706;
    reg [7:0] _708;
    wire [7:0] _709;
    wire [7:0] _710;
    wire [7:0] _711;
    reg [7:0] _702;
    wire [7:0] _703;
    wire [7:0] _704;
    reg [7:0] _712;
    wire [7:0] _27;
    reg [7:0] _175;
    wire [7:0] _719;
    reg [7:0] _721;
    wire [7:0] _722;
    wire [7:0] _723;
    wire [7:0] _724;
    reg [7:0] _715;
    wire [7:0] _716;
    wire [7:0] _717;
    reg [7:0] _725;
    wire [7:0] _28;
    reg [7:0] _173;
    wire [7:0] _732;
    reg [7:0] _734;
    wire [7:0] _735;
    wire [7:0] _736;
    wire [7:0] _737;
    reg [7:0] _728;
    wire [7:0] _729;
    wire [7:0] _730;
    reg [7:0] _738;
    wire [7:0] _29;
    reg [7:0] _171;
    wire [7:0] _745;
    reg [7:0] _747;
    wire [7:0] _748;
    wire [7:0] _749;
    wire [7:0] _750;
    reg [7:0] _741;
    wire [7:0] _742;
    wire [7:0] _743;
    reg [7:0] _751;
    wire [7:0] _30;
    reg [7:0] _169;
    wire [7:0] _758;
    reg [7:0] _760;
    wire [7:0] _761;
    wire [7:0] _762;
    wire [7:0] _763;
    reg [7:0] _754;
    wire [7:0] _755;
    wire [7:0] _756;
    reg [7:0] _764;
    wire [7:0] _31;
    reg [7:0] _167;
    wire [7:0] _771;
    reg [7:0] _773;
    wire [7:0] _774;
    wire [7:0] _775;
    wire [7:0] _776;
    reg [7:0] _767;
    wire [7:0] _768;
    wire [7:0] _769;
    reg [7:0] _777;
    wire [7:0] _32;
    reg [7:0] _165;
    wire [7:0] _785;
    reg [7:0] _787;
    wire [7:0] _788;
    wire [7:0] _789;
    wire [7:0] _790;
    reg [7:0] _781;
    wire [7:0] _782;
    wire [7:0] _783;
    reg [7:0] _791;
    wire [7:0] _33;
    reg [7:0] _163;
    wire [3:0] _793;
    wire [3:0] _794;
    wire [3:0] _795;
    wire [3:0] _796;
    wire [3:0] _797;
    reg [3:0] _798;
    wire [3:0] _34;
    reg [3:0] _225;
    wire [3:0] _1201;
    wire [3:0] _1198;
    wire [3:0] _1199;
    wire [2:0] _90;
    wire [2:0] _806;
    wire [2:0] _807;
    wire [2:0] _808;
    wire _193;
    wire [2:0] _800;
    wire [2:0] _801;
    wire [2:0] _802;
    wire [2:0] _803;
    reg [2:0] _809;
    wire [2:0] _35;
    reg [2:0] _235;
    wire _805;
    wire [2:0] _1194;
    wire [2:0] _1188;
    wire [2:0] _1190;
    wire [2:0] _130;
    wire [2:0] _822;
    reg [2:0] _824;
    reg [2:0] _819;
    reg [2:0] _815;
    wire [2:0] _816;
    wire [2:0] _820;
    wire [2:0] _825;
    reg [2:0] _811;
    wire [2:0] _812;
    wire [2:0] _813;
    reg [2:0] _826;
    wire [2:0] _36;
    reg [2:0] _128;
    wire [2:0] _839;
    reg [2:0] _841;
    reg [2:0] _836;
    reg [2:0] _832;
    wire [2:0] _833;
    wire [2:0] _837;
    wire [2:0] _842;
    reg [2:0] _828;
    wire [2:0] _829;
    wire [2:0] _830;
    reg [2:0] _843;
    wire [2:0] _37;
    reg [2:0] _126;
    wire [2:0] _856;
    reg [2:0] _858;
    reg [2:0] _853;
    reg [2:0] _849;
    wire [2:0] _850;
    wire [2:0] _854;
    wire [2:0] _859;
    reg [2:0] _845;
    wire [2:0] _846;
    wire [2:0] _847;
    reg [2:0] _860;
    wire [2:0] _38;
    reg [2:0] _124;
    wire [2:0] _873;
    reg [2:0] _875;
    reg [2:0] _870;
    reg [2:0] _866;
    wire [2:0] _867;
    wire [2:0] _871;
    wire [2:0] _876;
    reg [2:0] _862;
    wire [2:0] _863;
    wire [2:0] _864;
    reg [2:0] _877;
    wire [2:0] _39;
    reg [2:0] _122;
    wire [2:0] _890;
    reg [2:0] _892;
    reg [2:0] _887;
    reg [2:0] _883;
    wire [2:0] _884;
    wire [2:0] _888;
    wire [2:0] _893;
    reg [2:0] _879;
    wire [2:0] _880;
    wire [2:0] _881;
    reg [2:0] _894;
    wire [2:0] _40;
    reg [2:0] _120;
    wire [2:0] _907;
    reg [2:0] _909;
    reg [2:0] _904;
    reg [2:0] _900;
    wire [2:0] _901;
    wire [2:0] _905;
    wire [2:0] _910;
    reg [2:0] _896;
    wire [2:0] _897;
    wire [2:0] _898;
    reg [2:0] _911;
    wire [2:0] _41;
    reg [2:0] _118;
    wire [2:0] _924;
    reg [2:0] _926;
    reg [2:0] _921;
    reg [2:0] _917;
    wire [2:0] _918;
    wire [2:0] _922;
    wire [2:0] _927;
    reg [2:0] _913;
    wire [2:0] _914;
    wire [2:0] _915;
    reg [2:0] _928;
    wire [2:0] _42;
    reg [2:0] _116;
    wire [2:0] _941;
    reg [2:0] _943;
    reg [2:0] _938;
    reg [2:0] _934;
    wire [2:0] _935;
    wire [2:0] _939;
    wire [2:0] _944;
    reg [2:0] _930;
    wire [2:0] _931;
    wire [2:0] _932;
    reg [2:0] _945;
    wire [2:0] _43;
    reg [2:0] _114;
    wire [2:0] _958;
    reg [2:0] _960;
    reg [2:0] _955;
    reg [2:0] _951;
    wire [2:0] _952;
    wire [2:0] _956;
    wire [2:0] _961;
    reg [2:0] _947;
    wire [2:0] _948;
    wire [2:0] _949;
    reg [2:0] _962;
    wire [2:0] _44;
    reg [2:0] _112;
    wire [2:0] _975;
    reg [2:0] _977;
    reg [2:0] _972;
    reg [2:0] _968;
    wire [2:0] _969;
    wire [2:0] _973;
    wire [2:0] _978;
    reg [2:0] _964;
    wire [2:0] _965;
    wire [2:0] _966;
    reg [2:0] _979;
    wire [2:0] _45;
    reg [2:0] _110;
    wire [2:0] _992;
    reg [2:0] _994;
    reg [2:0] _989;
    reg [2:0] _985;
    wire [2:0] _986;
    wire [2:0] _990;
    wire [2:0] _995;
    reg [2:0] _981;
    wire [2:0] _982;
    wire [2:0] _983;
    reg [2:0] _996;
    wire [2:0] _46;
    reg [2:0] _108;
    wire [2:0] _1176;
    reg [2:0] _1178;
    reg [2:0] _1173;
    reg [2:0] _1170;
    wire [2:0] _1171;
    wire [7:0] _997;
    reg [7:0] _999;
    wire [7:0] _47;
    reg [7:0] _158;
    wire [7:0] _160;
    wire [7:0] _1008;
    reg [7:0] _1009;
    reg [7:0] _1005;
    wire [7:0] _1006;
    wire [7:0] _1010;
    wire [7:0] _1011;
    reg [7:0] _1001;
    wire [7:0] _1002;
    wire [7:0] _1003;
    reg [7:0] _1012;
    wire [7:0] _48;
    reg [7:0] _155;
    wire [7:0] _1021;
    reg [7:0] _1022;
    reg [7:0] _1018;
    wire [7:0] _1019;
    wire [7:0] _1023;
    wire [7:0] _1024;
    reg [7:0] _1014;
    wire [7:0] _1015;
    wire [7:0] _1016;
    reg [7:0] _1025;
    wire [7:0] _49;
    reg [7:0] _153;
    wire [7:0] _1034;
    reg [7:0] _1035;
    reg [7:0] _1031;
    wire [7:0] _1032;
    wire [7:0] _1036;
    wire [7:0] _1037;
    reg [7:0] _1027;
    wire [7:0] _1028;
    wire [7:0] _1029;
    reg [7:0] _1038;
    wire [7:0] _50;
    reg [7:0] _151;
    wire [7:0] _1047;
    reg [7:0] _1048;
    reg [7:0] _1044;
    wire [7:0] _1045;
    wire [7:0] _1049;
    wire [7:0] _1050;
    reg [7:0] _1040;
    wire [7:0] _1041;
    wire [7:0] _1042;
    reg [7:0] _1051;
    wire [7:0] _51;
    reg [7:0] _149;
    wire [7:0] _1060;
    reg [7:0] _1061;
    reg [7:0] _1057;
    wire [7:0] _1058;
    wire [7:0] _1062;
    wire [7:0] _1063;
    reg [7:0] _1053;
    wire [7:0] _1054;
    wire [7:0] _1055;
    reg [7:0] _1064;
    wire [7:0] _52;
    reg [7:0] _147;
    wire [7:0] _1073;
    reg [7:0] _1074;
    reg [7:0] _1070;
    wire [7:0] _1071;
    wire [7:0] _1075;
    wire [7:0] _1076;
    reg [7:0] _1066;
    wire [7:0] _1067;
    wire [7:0] _1068;
    reg [7:0] _1077;
    wire [7:0] _53;
    reg [7:0] _145;
    wire [7:0] _1086;
    reg [7:0] _1087;
    reg [7:0] _1083;
    wire [7:0] _1084;
    wire [7:0] _1088;
    wire [7:0] _1089;
    reg [7:0] _1079;
    wire [7:0] _1080;
    wire [7:0] _1081;
    reg [7:0] _1090;
    wire [7:0] _54;
    reg [7:0] _143;
    wire [7:0] _1099;
    reg [7:0] _1100;
    reg [7:0] _1096;
    wire [7:0] _1097;
    wire [7:0] _1101;
    wire [7:0] _1102;
    reg [7:0] _1092;
    wire [7:0] _1093;
    wire [7:0] _1094;
    reg [7:0] _1103;
    wire [7:0] _55;
    reg [7:0] _141;
    wire [7:0] _1112;
    reg [7:0] _1113;
    reg [7:0] _1109;
    wire [7:0] _1110;
    wire [7:0] _1114;
    wire [7:0] _1115;
    reg [7:0] _1105;
    wire [7:0] _1106;
    wire [7:0] _1107;
    reg [7:0] _1116;
    wire [7:0] _56;
    reg [7:0] _139;
    wire [7:0] _1125;
    reg [7:0] _1126;
    reg [7:0] _1122;
    wire [7:0] _1123;
    wire [7:0] _1127;
    wire [7:0] _1128;
    reg [7:0] _1118;
    wire [7:0] _1119;
    wire [7:0] _1120;
    reg [7:0] _1129;
    wire [7:0] _57;
    reg [7:0] _137;
    wire [7:0] _1138;
    reg [7:0] _1139;
    reg [7:0] _1135;
    wire [7:0] _1136;
    wire [7:0] _1140;
    wire [7:0] _1141;
    reg [7:0] _1131;
    wire [7:0] _1132;
    wire [7:0] _1133;
    reg [7:0] _1142;
    wire [7:0] _58;
    reg [7:0] _135;
    wire [7:0] _1158;
    reg [7:0] _1160;
    reg [7:0] _1155;
    wire [7:0] _1145;
    wire [7:0] _1146;
    reg [7:0] _1148;
    wire [7:0] _59;
    reg [7:0] _188;
    wire [7:0] _190;
    wire _191;
    wire [7:0] _1156;
    wire [7:0] _1161;
    wire [7:0] _1162;
    reg [7:0] _1151;
    wire [7:0] _1152;
    wire [7:0] _1153;
    reg [7:0] _1163;
    wire [7:0] _60;
    reg [7:0] _133;
    reg [7:0] _156;
    wire _161;
    wire [2:0] _1174;
    wire [2:0] _1179;
    wire [3:0] _634;
    reg [2:0] _1166;
    wire [2:0] _1167;
    wire [2:0] _1168;
    reg [2:0] _1180;
    wire [2:0] _61;
    reg [2:0] _106;
    reg [2:0] _129;
    wire _131;
    wire [2:0] _1192;
    wire [2:0] _1185;
    wire [3:0] _97;
    wire _98;
    wire [2:0] _1183;
    wire [2:0] _1186;
    reg [2:0] _1195;
    wire [2:0] _62;
    reg [2:0] _89;
    wire _91;
    wire [3:0] _1200;
    reg [3:0] _1202;
    wire [3:0] _63;
    reg [3:0] _93;
    reg [7:0] _186;
    wire [3:0] _221;
    wire _222;
    wire _219;
    wire [3:0] _216;
    wire _217;
    wire _220;
    wire _223;
    wire [7:0] _227;
    wire [7:0] _238;
    wire [3:0] _1205;
    reg [3:0] _1206;
    wire [3:0] _64;
    wire [15:0] _341;
    reg [15:0] _342;
    wire [15:0] _1318;
    wire _1320;
    wire _1321;
    wire _1352;
    wire _1355;
    wire [3:0] _1356;
    wire [3:0] _87;
    wire [3:0] _1313;
    wire [3:0] _1314;
    wire [3:0] _1312;
    wire [3:0] _1309;
    wire [2:0] _1303;
    wire [2:0] _1300;
    wire _1301;
    wire [2:0] _1304;
    wire [3:0] _1212;
    wire [3:0] _1213;
    wire [3:0] _1210;
    reg [3:0] _1214;
    wire [3:0] _65;
    reg [3:0] _95;
    wire _263;
    wire [7:0] _1222;
    reg [7:0] _1224;
    wire [7:0] _1225;
    reg [7:0] _1218;
    wire [7:0] _1219;
    wire [7:0] _1220;
    reg [7:0] _1226;
    wire [7:0] _66;
    reg [7:0] _257;
    wire [7:0] _1232;
    reg [7:0] _1234;
    wire [7:0] _1235;
    reg [7:0] _1228;
    wire [7:0] _1229;
    wire [7:0] _1230;
    reg [7:0] _1236;
    wire [7:0] _67;
    reg [7:0] _255;
    wire [7:0] _1242;
    reg [7:0] _1244;
    wire [7:0] _1245;
    reg [7:0] _1238;
    wire [7:0] _1239;
    wire [7:0] _1240;
    reg [7:0] _1246;
    wire [7:0] _68;
    reg [7:0] _253;
    wire [7:0] _1252;
    reg [7:0] _1254;
    wire [7:0] _1255;
    reg [7:0] _1248;
    wire [7:0] _1249;
    wire [7:0] _1250;
    reg [7:0] _1256;
    wire [7:0] _69;
    reg [7:0] _251;
    wire [7:0] _1262;
    reg [7:0] _1264;
    wire [7:0] _1265;
    reg [7:0] _1258;
    wire [7:0] _1259;
    wire [7:0] _1260;
    reg [7:0] _1266;
    wire [7:0] _70;
    reg [7:0] _249;
    wire [7:0] _1272;
    reg [7:0] _1274;
    wire [7:0] _1275;
    wire [7:0] _72;
    wire [2:0] _1215;
    wire [2:0] _1216;
    reg [7:0] _1268;
    wire [7:0] _1269;
    wire [7:0] _1270;
    reg [7:0] _1276;
    wire [7:0] _73;
    reg [7:0] _247;
    reg [7:0] _258;
    wire _260;
    wire _261;
    wire _264;
    wire [2:0] _1305;
    wire [3:0] _1207;
    wire _75;
    wire _77;
    wire [3:0] _1286;
    wire [3:0] _1287;
    wire [3:0] _1282;
    wire [3:0] _1283;
    wire [3:0] _1284;
    reg [3:0] _1288;
    wire [3:0] _78;
    reg [3:0] _1204;
    wire _1208;
    wire [2:0] _1299;
    wire _1144;
    wire [2:0] _1294;
    wire [2:0] _1292;
    wire _1280;
    wire [2:0] _1295;
    wire [2:0] _1296;
    wire [2:0] _1297;
    wire [2:0] _1290;
    reg [2:0] _1306;
    wire [2:0] _79;
    reg [2:0] _245;
    wire _1278;
    wire [3:0] _1310;
    wire [3:0] _1311;
    wire _81;
    wire [3:0] _1308;
    reg [3:0] _1365;
    wire [3:0] _82;
    (* fsm_encoding="one_hot" *)
    reg [3:0] _85;
    wire _1366;
    wire _1368;
    assign _99 = 1'b0;
    assign _194 = _193 ? vdd : _100;
    assign _195 = _191 ? _100 : _194;
    assign _196 = _161 ? _100 : _195;
    assign _197 = _131 ? _100 : _196;
    assign _102 = _98 ? vdd : _100;
    assign _103 = _91 ? _100 : _102;
    always @* begin
        case (_85)
        4'b0101:
            _199 <= gnd;
        4'b1001:
            _199 <= _103;
        4'b1010:
            _199 <= _197;
        default:
            _199 <= _100;
        endcase
    end
    assign _1 = _199;
    always @(posedge _77) begin
        if (_75)
            _100 <= _99;
        else
            _100 <= _1;
    end
    assign _204 = _193 ? gnd : _201;
    assign _205 = _191 ? _201 : _204;
    assign _206 = _161 ? _201 : _205;
    assign _207 = _131 ? _201 : _206;
    assign _202 = _98 ? vdd : _201;
    assign _203 = _91 ? _201 : _202;
    always @* begin
        case (_85)
        4'b0101:
            _208 <= gnd;
        4'b1001:
            _208 <= _203;
        4'b1010:
            _208 <= _207;
        default:
            _208 <= _201;
        endcase
    end
    assign _2 = _208;
    always @(posedge _77) begin
        if (_75)
            _201 <= _99;
        else
            _201 <= _2;
    end
    assign _210 = _201 & _100;
    assign _209 = 7'b0000000;
    assign _211 = { _209,
                    _210 };
    assign _213 = _212 == _85;
    assign _214 = _212 == _85;
    assign _1367 = _604 == _85;
    assign _84 = 4'b0000;
    assign _7 = m_tready;
    assign _1364 = _7 ? _527 : _85;
    assign _1363 = _805 ? _216 : _198;
    assign _1359 = _193 ? _212 : _216;
    assign _1360 = _191 ? _602 : _1359;
    assign _1361 = _161 ? _602 : _1360;
    assign _1362 = _131 ? _602 : _1361;
    assign _212 = 4'b1110;
    assign _1357 = _98 ? _212 : _602;
    assign _1358 = _91 ? _602 : _1357;
    assign _198 = 4'b1010;
    assign _104 = 4'b1001;
    assign _1353 = _238 < _188;
    assign _1354 = ~ _1353;
    assign _1349 = 16'b0000000000000000;
    assign _1345 = 16'b0000000000000001;
    assign _1340 = 8'b00000000;
    assign _1339 = _1338[7:0];
    assign _1341 = { _1339,
                     _1340 };
    assign _1335 = _1334[11:0];
    assign _1337 = { _1335,
                     _84 };
    assign _1332 = 2'b00;
    assign _1331 = _1330[13:0];
    assign _1333 = { _1331,
                     _1332 };
    assign _1329 = 16'b0000000000000010;
    assign _1327 = _1322[0:0];
    assign _1330 = _1327 ? _1329 : _1345;
    assign _1326 = _1322[1:1];
    assign _1334 = _1326 ? _1333 : _1330;
    assign _1325 = _1322[2:2];
    assign _1338 = _1325 ? _1337 : _1334;
    assign _1324 = _1322[3:3];
    assign _1342 = _1324 ? _1341 : _1338;
    assign _1322 = _158[4:0];
    assign _1323 = _1322[4:4];
    assign _1344 = _1323 ? _1349 : _1342;
    assign _1346 = _1344 - _1345;
    assign _1347 = ~ _1346;
    assign _1348 = _626 & _1347;
    assign _1350 = _1348 == _1349;
    assign _1351 = ~ _1350;
    assign _242 = _241 ? vdd : gnd;
    assign gnd = 1'b0;
    assign _240 = _239 ? vdd : gnd;
    assign vdd = 1'b1;
    always @* begin
        case (_85)
        4'b0011:
            _243 <= vdd;
        4'b1001:
            _243 <= _240;
        4'b1101:
            _243 <= _242;
        default:
            _243 <= gnd;
        endcase
    end
    assign _8 = _243;
    assign _629 = ~ _626;
    assign _630 = _342 & _629;
    assign _241 = _238 < _188;
    assign _631 = _241 ? _630 : _1349;
    assign _623 = _622[7:0];
    assign _625 = { _623,
                    _1340 };
    assign _619 = _618[11:0];
    assign _621 = { _619,
                    _84 };
    assign _615 = _614[13:0];
    assign _617 = { _615,
                    _1332 };
    assign _611 = _610[14:0];
    assign _613 = { _611,
                    _99 };
    assign _604 = 4'b0010;
    assign _602 = 4'b0110;
    always @* begin
        case (_361)
        0:
            _606 <= _602;
        1:
            _606 <= _212;
        2:
            _606 <= _604;
        default:
            _606 <= _84;
        endcase
    end
    assign _598 = 4'b0111;
    assign _597 = 4'b0100;
    always @* begin
        case (_361)
        0:
            _601 <= _597;
        1:
            _601 <= _598;
        2:
            _601 <= _602;
        default:
            _601 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _596 <= _84;
        1:
            _596 <= _212;
        2:
            _596 <= _597;
        default:
            _596 <= _212;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _591 <= _212;
        1:
            _591 <= _597;
        2:
            _591 <= _212;
        default:
            _591 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _586 <= _602;
        1:
            _586 <= _212;
        2:
            _586 <= _604;
        default:
            _586 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _581 <= _84;
        1:
            _581 <= _212;
        2:
            _581 <= _597;
        default:
            _581 <= _212;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _576 <= _597;
        1:
            _576 <= _598;
        2:
            _576 <= _602;
        default:
            _576 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _571 <= _598;
        1:
            _571 <= _604;
        2:
            _571 <= _598;
        default:
            _571 <= _84;
        endcase
    end
    always @* begin
        case (_360)
        0:
            _607 <= _571;
        1:
            _607 <= _576;
        2:
            _607 <= _581;
        3:
            _607 <= _586;
        4:
            _607 <= _591;
        5:
            _607 <= _596;
        6:
            _607 <= _601;
        default:
            _607 <= _606;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _565 <= _597;
        1:
            _565 <= _212;
        2:
            _565 <= _602;
        default:
            _565 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _560 <= _602;
        1:
            _560 <= _598;
        2:
            _560 <= _604;
        default:
            _560 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _555 <= _84;
        1:
            _555 <= _212;
        2:
            _555 <= _597;
        default:
            _555 <= _212;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _550 <= _212;
        1:
            _550 <= _597;
        2:
            _550 <= _212;
        default:
            _550 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _545 <= _597;
        1:
            _545 <= _212;
        2:
            _545 <= _602;
        default:
            _545 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _540 <= _84;
        1:
            _540 <= _212;
        2:
            _540 <= _597;
        default:
            _540 <= _212;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _535 <= _602;
        1:
            _535 <= _598;
        2:
            _535 <= _604;
        default:
            _535 <= _84;
        endcase
    end
    assign _527 = 4'b0001;
    always @* begin
        case (_361)
        0:
            _530 <= _598;
        1:
            _530 <= _527;
        2:
            _530 <= _598;
        default:
            _530 <= _84;
        endcase
    end
    always @* begin
        case (_360)
        0:
            _566 <= _530;
        1:
            _566 <= _535;
        2:
            _566 <= _540;
        3:
            _566 <= _545;
        4:
            _566 <= _550;
        5:
            _566 <= _555;
        6:
            _566 <= _560;
        default:
            _566 <= _565;
        endcase
    end
    assign _521 = 4'b1100;
    always @* begin
        case (_361)
        0:
            _524 <= _602;
        1:
            _524 <= _521;
        2:
            _524 <= _602;
        default:
            _524 <= _84;
        endcase
    end
    assign _516 = 4'b0011;
    always @* begin
        case (_361)
        0:
            _519 <= _602;
        1:
            _519 <= _516;
        2:
            _519 <= _602;
        default:
            _519 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _514 <= _602;
        1:
            _514 <= _516;
        2:
            _514 <= _602;
        default:
            _514 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _509 <= _602;
        1:
            _509 <= _521;
        2:
            _509 <= _602;
        default:
            _509 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _504 <= _602;
        1:
            _504 <= _598;
        2:
            _504 <= _602;
        default:
            _504 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _499 <= _602;
        1:
            _499 <= _598;
        2:
            _499 <= _602;
        default:
            _499 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _494 <= _602;
        1:
            _494 <= _598;
        2:
            _494 <= _602;
        default:
            _494 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _489 <= _602;
        1:
            _489 <= _598;
        2:
            _489 <= _602;
        default:
            _489 <= _84;
        endcase
    end
    always @* begin
        case (_360)
        0:
            _525 <= _489;
        1:
            _525 <= _494;
        2:
            _525 <= _499;
        3:
            _525 <= _504;
        4:
            _525 <= _509;
        5:
            _525 <= _514;
        6:
            _525 <= _519;
        default:
            _525 <= _524;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _483 <= _521;
        1:
            _483 <= _602;
        2:
            _483 <= _602;
        default:
            _483 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _478 <= _602;
        1:
            _478 <= _598;
        2:
            _478 <= _516;
        default:
            _478 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _473 <= _84;
        1:
            _473 <= _602;
        2:
            _473 <= _212;
        default:
            _473 <= _516;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _468 <= _521;
        1:
            _468 <= _212;
        2:
            _468 <= _602;
        default:
            _468 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _463 <= _602;
        1:
            _463 <= _602;
        2:
            _463 <= _516;
        default:
            _463 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _458 <= _84;
        1:
            _458 <= _521;
        2:
            _458 <= _212;
        default:
            _458 <= _602;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _453 <= _521;
        1:
            _453 <= _602;
        2:
            _453 <= _602;
        default:
            _453 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _448 <= _602;
        1:
            _448 <= _598;
        2:
            _448 <= _516;
        default:
            _448 <= _84;
        endcase
    end
    always @* begin
        case (_360)
        0:
            _484 <= _448;
        1:
            _484 <= _453;
        2:
            _484 <= _458;
        3:
            _484 <= _463;
        4:
            _484 <= _468;
        5:
            _484 <= _473;
        6:
            _484 <= _478;
        default:
            _484 <= _483;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _442 <= _604;
        1:
            _442 <= _212;
        2:
            _442 <= _602;
        default:
            _442 <= _84;
        endcase
    end
    assign _436 = 4'b1000;
    always @* begin
        case (_361)
        0:
            _437 <= _84;
        1:
            _437 <= _521;
        2:
            _437 <= _602;
        default:
            _437 <= _436;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _432 <= _84;
        1:
            _432 <= _212;
        2:
            _432 <= _602;
        default:
            _432 <= _516;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _427 <= _521;
        1:
            _427 <= _212;
        2:
            _427 <= _602;
        default:
            _427 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _422 <= _436;
        1:
            _422 <= _212;
        2:
            _422 <= _602;
        default:
            _422 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _417 <= _84;
        1:
            _417 <= _212;
        2:
            _417 <= _602;
        default:
            _417 <= _521;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _412 <= _602;
        1:
            _412 <= _598;
        2:
            _412 <= _527;
        default:
            _412 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _407 <= _516;
        1:
            _407 <= _602;
        2:
            _407 <= _598;
        default:
            _407 <= _84;
        endcase
    end
    always @* begin
        case (_360)
        0:
            _443 <= _407;
        1:
            _443 <= _412;
        2:
            _443 <= _417;
        3:
            _443 <= _422;
        4:
            _443 <= _427;
        5:
            _443 <= _432;
        6:
            _443 <= _437;
        default:
            _443 <= _442;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _401 <= _436;
        1:
            _401 <= _212;
        2:
            _401 <= _602;
        default:
            _401 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _396 <= _84;
        1:
            _396 <= _598;
        2:
            _396 <= _602;
        default:
            _396 <= _597;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _391 <= _84;
        1:
            _391 <= _516;
        2:
            _391 <= _602;
        default:
            _391 <= _521;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _386 <= _602;
        1:
            _386 <= _521;
        2:
            _386 <= _602;
        default:
            _386 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _381 <= _521;
        1:
            _381 <= _212;
        2:
            _381 <= _602;
        default:
            _381 <= _84;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _376 <= _84;
        1:
            _376 <= _212;
        2:
            _376 <= _602;
        default:
            _376 <= _602;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _371 <= _602;
        1:
            _371 <= _598;
        2:
            _371 <= _516;
        default:
            _371 <= _84;
        endcase
    end
    assign _361 = _236[1:0];
    always @* begin
        case (_361)
        0:
            _366 <= _602;
        1:
            _366 <= _602;
        2:
            _366 <= _598;
        default:
            _366 <= _84;
        endcase
    end
    always @* begin
        case (_225)
        0:
            _359 <= _106;
        1:
            _359 <= _108;
        2:
            _359 <= _110;
        3:
            _359 <= _112;
        4:
            _359 <= _114;
        5:
            _359 <= _116;
        6:
            _359 <= _118;
        7:
            _359 <= _120;
        8:
            _359 <= _122;
        9:
            _359 <= _124;
        10:
            _359 <= _126;
        default:
            _359 <= _128;
        endcase
    end
    assign _360 = _223 ? _359 : _129;
    always @* begin
        case (_360)
        0:
            _402 <= _366;
        1:
            _402 <= _371;
        2:
            _402 <= _376;
        3:
            _402 <= _381;
        4:
            _402 <= _386;
        5:
            _402 <= _391;
        6:
            _402 <= _396;
        default:
            _402 <= _401;
        endcase
    end
    always @* begin
        case (_225)
        0:
            _357 <= _333;
        1:
            _357 <= _327;
        2:
            _357 <= _321;
        3:
            _357 <= _315;
        4:
            _357 <= _309;
        5:
            _357 <= _303;
        6:
            _357 <= _297;
        7:
            _357 <= _291;
        8:
            _357 <= _285;
        9:
            _357 <= _279;
        10:
            _357 <= _273;
        default:
            _357 <= _266;
        endcase
    end
    assign _265 = 3'b000;
    always @* begin
        case (_95)
        4'b1011:
            _268 <= _245;
        default:
            _268 <= _266;
        endcase
    end
    assign _269 = _264 ? _268 : _266;
    always @* begin
        case (_85)
        4'b0100:
            _271 <= _269;
        default:
            _271 <= _266;
        endcase
    end
    assign _9 = _271;
    always @(posedge _77) begin
        if (_75)
            _266 <= _265;
        else
            _266 <= _9;
    end
    always @* begin
        case (_95)
        4'b1010:
            _275 <= _245;
        default:
            _275 <= _273;
        endcase
    end
    assign _276 = _264 ? _275 : _273;
    always @* begin
        case (_85)
        4'b0100:
            _277 <= _276;
        default:
            _277 <= _273;
        endcase
    end
    assign _10 = _277;
    always @(posedge _77) begin
        if (_75)
            _273 <= _265;
        else
            _273 <= _10;
    end
    always @* begin
        case (_95)
        4'b1001:
            _281 <= _245;
        default:
            _281 <= _279;
        endcase
    end
    assign _282 = _264 ? _281 : _279;
    always @* begin
        case (_85)
        4'b0100:
            _283 <= _282;
        default:
            _283 <= _279;
        endcase
    end
    assign _11 = _283;
    always @(posedge _77) begin
        if (_75)
            _279 <= _265;
        else
            _279 <= _11;
    end
    always @* begin
        case (_95)
        4'b1000:
            _287 <= _245;
        default:
            _287 <= _285;
        endcase
    end
    assign _288 = _264 ? _287 : _285;
    always @* begin
        case (_85)
        4'b0100:
            _289 <= _288;
        default:
            _289 <= _285;
        endcase
    end
    assign _12 = _289;
    always @(posedge _77) begin
        if (_75)
            _285 <= _265;
        else
            _285 <= _12;
    end
    always @* begin
        case (_95)
        4'b0111:
            _293 <= _245;
        default:
            _293 <= _291;
        endcase
    end
    assign _294 = _264 ? _293 : _291;
    always @* begin
        case (_85)
        4'b0100:
            _295 <= _294;
        default:
            _295 <= _291;
        endcase
    end
    assign _13 = _295;
    always @(posedge _77) begin
        if (_75)
            _291 <= _265;
        else
            _291 <= _13;
    end
    always @* begin
        case (_95)
        4'b0110:
            _299 <= _245;
        default:
            _299 <= _297;
        endcase
    end
    assign _300 = _264 ? _299 : _297;
    always @* begin
        case (_85)
        4'b0100:
            _301 <= _300;
        default:
            _301 <= _297;
        endcase
    end
    assign _14 = _301;
    always @(posedge _77) begin
        if (_75)
            _297 <= _265;
        else
            _297 <= _14;
    end
    always @* begin
        case (_95)
        4'b0101:
            _305 <= _245;
        default:
            _305 <= _303;
        endcase
    end
    assign _306 = _264 ? _305 : _303;
    always @* begin
        case (_85)
        4'b0100:
            _307 <= _306;
        default:
            _307 <= _303;
        endcase
    end
    assign _15 = _307;
    always @(posedge _77) begin
        if (_75)
            _303 <= _265;
        else
            _303 <= _15;
    end
    always @* begin
        case (_95)
        4'b0100:
            _311 <= _245;
        default:
            _311 <= _309;
        endcase
    end
    assign _312 = _264 ? _311 : _309;
    always @* begin
        case (_85)
        4'b0100:
            _313 <= _312;
        default:
            _313 <= _309;
        endcase
    end
    assign _16 = _313;
    always @(posedge _77) begin
        if (_75)
            _309 <= _265;
        else
            _309 <= _16;
    end
    always @* begin
        case (_95)
        4'b0011:
            _317 <= _245;
        default:
            _317 <= _315;
        endcase
    end
    assign _318 = _264 ? _317 : _315;
    always @* begin
        case (_85)
        4'b0100:
            _319 <= _318;
        default:
            _319 <= _315;
        endcase
    end
    assign _17 = _319;
    always @(posedge _77) begin
        if (_75)
            _315 <= _265;
        else
            _315 <= _17;
    end
    always @* begin
        case (_95)
        4'b0010:
            _323 <= _245;
        default:
            _323 <= _321;
        endcase
    end
    assign _324 = _264 ? _323 : _321;
    always @* begin
        case (_85)
        4'b0100:
            _325 <= _324;
        default:
            _325 <= _321;
        endcase
    end
    assign _18 = _325;
    always @(posedge _77) begin
        if (_75)
            _321 <= _265;
        else
            _321 <= _18;
    end
    always @* begin
        case (_95)
        4'b0001:
            _329 <= _245;
        default:
            _329 <= _327;
        endcase
    end
    assign _330 = _264 ? _329 : _327;
    always @* begin
        case (_85)
        4'b0100:
            _331 <= _330;
        default:
            _331 <= _327;
        endcase
    end
    assign _19 = _331;
    always @(posedge _77) begin
        if (_75)
            _327 <= _265;
        else
            _327 <= _19;
    end
    always @* begin
        case (_95)
        4'b0000:
            _335 <= _245;
        default:
            _335 <= _333;
        endcase
    end
    assign _336 = _264 ? _335 : _333;
    always @* begin
        case (_85)
        4'b0100:
            _337 <= _336;
        default:
            _337 <= _333;
        endcase
    end
    assign _20 = _337;
    always @(posedge _77) begin
        if (_75)
            _333 <= _265;
        else
            _333 <= _20;
    end
    always @* begin
        case (_93)
        0:
            _356 <= _333;
        1:
            _356 <= _327;
        2:
            _356 <= _321;
        3:
            _356 <= _315;
        4:
            _356 <= _309;
        5:
            _356 <= _303;
        6:
            _356 <= _297;
        7:
            _356 <= _291;
        8:
            _356 <= _285;
        9:
            _356 <= _279;
        10:
            _356 <= _273;
        default:
            _356 <= _266;
        endcase
    end
    assign _358 = _223 ? _357 : _356;
    always @* begin
        case (_358)
        0:
            _608 <= _402;
        1:
            _608 <= _443;
        2:
            _608 <= _484;
        3:
            _608 <= _525;
        4:
            _608 <= _566;
        default:
            _608 <= _607;
        endcase
    end
    assign _355 = 12'b000000000000;
    assign _609 = { _355,
                    _608 };
    assign _352 = _238 < _188;
    assign _350 = 3'b100;
    assign _351 = _236 < _350;
    assign _353 = _351 & _352;
    assign _610 = _353 ? _609 : _1349;
    assign _349 = _345[0:0];
    assign _614 = _349 ? _613 : _610;
    assign _348 = _345[1:1];
    assign _618 = _348 ? _617 : _614;
    assign _347 = _345[2:2];
    assign _622 = _347 ? _621 : _618;
    always @* begin
        case (_225)
        0:
            _343 <= _133;
        1:
            _343 <= _135;
        2:
            _343 <= _137;
        3:
            _343 <= _139;
        4:
            _343 <= _141;
        5:
            _343 <= _143;
        6:
            _343 <= _145;
        7:
            _343 <= _147;
        8:
            _343 <= _149;
        9:
            _343 <= _151;
        10:
            _343 <= _153;
        default:
            _343 <= _155;
        endcase
    end
    assign _344 = _223 ? _343 : _156;
    assign _345 = _344[3:0];
    assign _346 = _345[3:3];
    assign _626 = _346 ? _625 : _622;
    assign _627 = _342 | _626;
    assign _239 = _238 < _188;
    assign _628 = _239 ? _627 : _1349;
    always @* begin
        case (_85)
        4'b0011:
            _632 <= _1349;
        4'b1001:
            _632 <= _628;
        4'b1101:
            _632 <= _631;
        default:
            _632 <= _1349;
        endcase
    end
    assign _21 = _632;
    always @(posedge _77) begin
        if (_8)
            _340[_64] <= _21;
    end
    assign _232 = _221 == _85;
    assign _230 = _521 == _85;
    assign _229 = _216 == _85;
    assign _231 = _229 | _230;
    assign _233 = _231 | _232;
    assign _236 = _233 ? _235 : _89;
    assign _228 = 5'b00000;
    assign _237 = { _228,
                    _236 };
    always @* begin
        case (_225)
        0:
            _226 <= _163;
        1:
            _226 <= _165;
        2:
            _226 <= _167;
        3:
            _226 <= _169;
        4:
            _226 <= _171;
        5:
            _226 <= _173;
        6:
            _226 <= _175;
        7:
            _226 <= _177;
        8:
            _226 <= _179;
        9:
            _226 <= _181;
        10:
            _226 <= _183;
        default:
            _226 <= _185;
        endcase
    end
    assign _640 = 8'b00000001;
    assign _641 = _185 + _640;
    always @* begin
        case (_93)
        4'b1011:
            _643 <= _641;
        default:
            _643 <= _185;
        endcase
    end
    assign _644 = _191 ? _643 : _185;
    assign _645 = _161 ? _185 : _644;
    assign _646 = _131 ? _185 : _645;
    always @* begin
        case (_634)
        4'b1011:
            _637 <= _1340;
        default:
            _637 <= _185;
        endcase
    end
    assign _638 = _98 ? _185 : _637;
    assign _639 = _91 ? _185 : _638;
    always @* begin
        case (_85)
        4'b1001:
            _647 <= _639;
        4'b1010:
            _647 <= _646;
        default:
            _647 <= _185;
        endcase
    end
    assign _22 = _647;
    always @(posedge _77) begin
        if (_75)
            _185 <= _1340;
        else
            _185 <= _22;
    end
    assign _654 = _183 + _640;
    always @* begin
        case (_93)
        4'b1010:
            _656 <= _654;
        default:
            _656 <= _183;
        endcase
    end
    assign _657 = _191 ? _656 : _183;
    assign _658 = _161 ? _183 : _657;
    assign _659 = _131 ? _183 : _658;
    always @* begin
        case (_634)
        4'b1010:
            _650 <= _1340;
        default:
            _650 <= _183;
        endcase
    end
    assign _651 = _98 ? _183 : _650;
    assign _652 = _91 ? _183 : _651;
    always @* begin
        case (_85)
        4'b1001:
            _660 <= _652;
        4'b1010:
            _660 <= _659;
        default:
            _660 <= _183;
        endcase
    end
    assign _23 = _660;
    always @(posedge _77) begin
        if (_75)
            _183 <= _1340;
        else
            _183 <= _23;
    end
    assign _667 = _181 + _640;
    always @* begin
        case (_93)
        4'b1001:
            _669 <= _667;
        default:
            _669 <= _181;
        endcase
    end
    assign _670 = _191 ? _669 : _181;
    assign _671 = _161 ? _181 : _670;
    assign _672 = _131 ? _181 : _671;
    always @* begin
        case (_634)
        4'b1001:
            _663 <= _1340;
        default:
            _663 <= _181;
        endcase
    end
    assign _664 = _98 ? _181 : _663;
    assign _665 = _91 ? _181 : _664;
    always @* begin
        case (_85)
        4'b1001:
            _673 <= _665;
        4'b1010:
            _673 <= _672;
        default:
            _673 <= _181;
        endcase
    end
    assign _24 = _673;
    always @(posedge _77) begin
        if (_75)
            _181 <= _1340;
        else
            _181 <= _24;
    end
    assign _680 = _179 + _640;
    always @* begin
        case (_93)
        4'b1000:
            _682 <= _680;
        default:
            _682 <= _179;
        endcase
    end
    assign _683 = _191 ? _682 : _179;
    assign _684 = _161 ? _179 : _683;
    assign _685 = _131 ? _179 : _684;
    always @* begin
        case (_634)
        4'b1000:
            _676 <= _1340;
        default:
            _676 <= _179;
        endcase
    end
    assign _677 = _98 ? _179 : _676;
    assign _678 = _91 ? _179 : _677;
    always @* begin
        case (_85)
        4'b1001:
            _686 <= _678;
        4'b1010:
            _686 <= _685;
        default:
            _686 <= _179;
        endcase
    end
    assign _25 = _686;
    always @(posedge _77) begin
        if (_75)
            _179 <= _1340;
        else
            _179 <= _25;
    end
    assign _693 = _177 + _640;
    always @* begin
        case (_93)
        4'b0111:
            _695 <= _693;
        default:
            _695 <= _177;
        endcase
    end
    assign _696 = _191 ? _695 : _177;
    assign _697 = _161 ? _177 : _696;
    assign _698 = _131 ? _177 : _697;
    always @* begin
        case (_634)
        4'b0111:
            _689 <= _1340;
        default:
            _689 <= _177;
        endcase
    end
    assign _690 = _98 ? _177 : _689;
    assign _691 = _91 ? _177 : _690;
    always @* begin
        case (_85)
        4'b1001:
            _699 <= _691;
        4'b1010:
            _699 <= _698;
        default:
            _699 <= _177;
        endcase
    end
    assign _26 = _699;
    always @(posedge _77) begin
        if (_75)
            _177 <= _1340;
        else
            _177 <= _26;
    end
    assign _706 = _175 + _640;
    always @* begin
        case (_93)
        4'b0110:
            _708 <= _706;
        default:
            _708 <= _175;
        endcase
    end
    assign _709 = _191 ? _708 : _175;
    assign _710 = _161 ? _175 : _709;
    assign _711 = _131 ? _175 : _710;
    always @* begin
        case (_634)
        4'b0110:
            _702 <= _1340;
        default:
            _702 <= _175;
        endcase
    end
    assign _703 = _98 ? _175 : _702;
    assign _704 = _91 ? _175 : _703;
    always @* begin
        case (_85)
        4'b1001:
            _712 <= _704;
        4'b1010:
            _712 <= _711;
        default:
            _712 <= _175;
        endcase
    end
    assign _27 = _712;
    always @(posedge _77) begin
        if (_75)
            _175 <= _1340;
        else
            _175 <= _27;
    end
    assign _719 = _173 + _640;
    always @* begin
        case (_93)
        4'b0101:
            _721 <= _719;
        default:
            _721 <= _173;
        endcase
    end
    assign _722 = _191 ? _721 : _173;
    assign _723 = _161 ? _173 : _722;
    assign _724 = _131 ? _173 : _723;
    always @* begin
        case (_634)
        4'b0101:
            _715 <= _1340;
        default:
            _715 <= _173;
        endcase
    end
    assign _716 = _98 ? _173 : _715;
    assign _717 = _91 ? _173 : _716;
    always @* begin
        case (_85)
        4'b1001:
            _725 <= _717;
        4'b1010:
            _725 <= _724;
        default:
            _725 <= _173;
        endcase
    end
    assign _28 = _725;
    always @(posedge _77) begin
        if (_75)
            _173 <= _1340;
        else
            _173 <= _28;
    end
    assign _732 = _171 + _640;
    always @* begin
        case (_93)
        4'b0100:
            _734 <= _732;
        default:
            _734 <= _171;
        endcase
    end
    assign _735 = _191 ? _734 : _171;
    assign _736 = _161 ? _171 : _735;
    assign _737 = _131 ? _171 : _736;
    always @* begin
        case (_634)
        4'b0100:
            _728 <= _1340;
        default:
            _728 <= _171;
        endcase
    end
    assign _729 = _98 ? _171 : _728;
    assign _730 = _91 ? _171 : _729;
    always @* begin
        case (_85)
        4'b1001:
            _738 <= _730;
        4'b1010:
            _738 <= _737;
        default:
            _738 <= _171;
        endcase
    end
    assign _29 = _738;
    always @(posedge _77) begin
        if (_75)
            _171 <= _1340;
        else
            _171 <= _29;
    end
    assign _745 = _169 + _640;
    always @* begin
        case (_93)
        4'b0011:
            _747 <= _745;
        default:
            _747 <= _169;
        endcase
    end
    assign _748 = _191 ? _747 : _169;
    assign _749 = _161 ? _169 : _748;
    assign _750 = _131 ? _169 : _749;
    always @* begin
        case (_634)
        4'b0011:
            _741 <= _1340;
        default:
            _741 <= _169;
        endcase
    end
    assign _742 = _98 ? _169 : _741;
    assign _743 = _91 ? _169 : _742;
    always @* begin
        case (_85)
        4'b1001:
            _751 <= _743;
        4'b1010:
            _751 <= _750;
        default:
            _751 <= _169;
        endcase
    end
    assign _30 = _751;
    always @(posedge _77) begin
        if (_75)
            _169 <= _1340;
        else
            _169 <= _30;
    end
    assign _758 = _167 + _640;
    always @* begin
        case (_93)
        4'b0010:
            _760 <= _758;
        default:
            _760 <= _167;
        endcase
    end
    assign _761 = _191 ? _760 : _167;
    assign _762 = _161 ? _167 : _761;
    assign _763 = _131 ? _167 : _762;
    always @* begin
        case (_634)
        4'b0010:
            _754 <= _1340;
        default:
            _754 <= _167;
        endcase
    end
    assign _755 = _98 ? _167 : _754;
    assign _756 = _91 ? _167 : _755;
    always @* begin
        case (_85)
        4'b1001:
            _764 <= _756;
        4'b1010:
            _764 <= _763;
        default:
            _764 <= _167;
        endcase
    end
    assign _31 = _764;
    always @(posedge _77) begin
        if (_75)
            _167 <= _1340;
        else
            _167 <= _31;
    end
    assign _771 = _165 + _640;
    always @* begin
        case (_93)
        4'b0001:
            _773 <= _771;
        default:
            _773 <= _165;
        endcase
    end
    assign _774 = _191 ? _773 : _165;
    assign _775 = _161 ? _165 : _774;
    assign _776 = _131 ? _165 : _775;
    always @* begin
        case (_634)
        4'b0001:
            _767 <= _1340;
        default:
            _767 <= _165;
        endcase
    end
    assign _768 = _98 ? _165 : _767;
    assign _769 = _91 ? _165 : _768;
    always @* begin
        case (_85)
        4'b1001:
            _777 <= _769;
        4'b1010:
            _777 <= _776;
        default:
            _777 <= _165;
        endcase
    end
    assign _32 = _777;
    always @(posedge _77) begin
        if (_75)
            _165 <= _1340;
        else
            _165 <= _32;
    end
    assign _785 = _163 + _640;
    always @* begin
        case (_93)
        4'b0000:
            _787 <= _785;
        default:
            _787 <= _163;
        endcase
    end
    assign _788 = _191 ? _787 : _163;
    assign _789 = _161 ? _163 : _788;
    assign _790 = _131 ? _163 : _789;
    always @* begin
        case (_634)
        4'b0000:
            _781 <= _1340;
        default:
            _781 <= _163;
        endcase
    end
    assign _782 = _98 ? _163 : _781;
    assign _783 = _91 ? _163 : _782;
    always @* begin
        case (_85)
        4'b0101:
            _791 <= _1340;
        4'b1001:
            _791 <= _783;
        4'b1010:
            _791 <= _790;
        default:
            _791 <= _163;
        endcase
    end
    assign _33 = _791;
    always @(posedge _77) begin
        if (_75)
            _163 <= _1340;
        else
            _163 <= _33;
    end
    assign _793 = _93 - _527;
    assign _794 = _193 ? _225 : _793;
    assign _795 = _191 ? _225 : _794;
    assign _796 = _161 ? _225 : _795;
    assign _797 = _131 ? _225 : _796;
    always @* begin
        case (_85)
        4'b1010:
            _798 <= _797;
        default:
            _798 <= _225;
        endcase
    end
    assign _34 = _798;
    always @(posedge _77) begin
        if (_75)
            _225 <= _84;
        else
            _225 <= _34;
    end
    assign _1201 = _805 ? _93 : _225;
    assign _1198 = _93 + _527;
    assign _1199 = _98 ? _93 : _1198;
    assign _90 = 3'b011;
    assign _806 = 3'b001;
    assign _807 = _235 + _806;
    assign _808 = _805 ? _807 : _235;
    assign _193 = _93 == _84;
    assign _800 = _193 ? _235 : _265;
    assign _801 = _191 ? _235 : _800;
    assign _802 = _161 ? _235 : _801;
    assign _803 = _131 ? _235 : _802;
    always @* begin
        case (_85)
        4'b1010:
            _809 <= _803;
        4'b1101:
            _809 <= _808;
        default:
            _809 <= _235;
        endcase
    end
    assign _35 = _809;
    always @(posedge _77) begin
        if (_75)
            _235 <= _265;
        else
            _235 <= _35;
    end
    assign _805 = _235 < _90;
    assign _1194 = _805 ? _89 : _265;
    assign _1188 = _191 ? _265 : _89;
    assign _1190 = _161 ? _265 : _1188;
    assign _130 = 3'b111;
    assign _822 = _128 + _806;
    always @* begin
        case (_93)
        4'b1011:
            _824 <= _822;
        default:
            _824 <= _128;
        endcase
    end
    always @* begin
        case (_93)
        4'b1011:
            _819 <= _265;
        default:
            _819 <= _128;
        endcase
    end
    always @* begin
        case (_93)
        4'b1011:
            _815 <= _265;
        default:
            _815 <= _128;
        endcase
    end
    assign _816 = _191 ? _815 : _128;
    assign _820 = _161 ? _819 : _816;
    assign _825 = _131 ? _824 : _820;
    always @* begin
        case (_634)
        4'b1011:
            _811 <= _265;
        default:
            _811 <= _128;
        endcase
    end
    assign _812 = _98 ? _128 : _811;
    assign _813 = _91 ? _128 : _812;
    always @* begin
        case (_85)
        4'b1001:
            _826 <= _813;
        4'b1010:
            _826 <= _825;
        default:
            _826 <= _128;
        endcase
    end
    assign _36 = _826;
    always @(posedge _77) begin
        if (_75)
            _128 <= _265;
        else
            _128 <= _36;
    end
    assign _839 = _126 + _806;
    always @* begin
        case (_93)
        4'b1010:
            _841 <= _839;
        default:
            _841 <= _126;
        endcase
    end
    always @* begin
        case (_93)
        4'b1010:
            _836 <= _265;
        default:
            _836 <= _126;
        endcase
    end
    always @* begin
        case (_93)
        4'b1010:
            _832 <= _265;
        default:
            _832 <= _126;
        endcase
    end
    assign _833 = _191 ? _832 : _126;
    assign _837 = _161 ? _836 : _833;
    assign _842 = _131 ? _841 : _837;
    always @* begin
        case (_634)
        4'b1010:
            _828 <= _265;
        default:
            _828 <= _126;
        endcase
    end
    assign _829 = _98 ? _126 : _828;
    assign _830 = _91 ? _126 : _829;
    always @* begin
        case (_85)
        4'b1001:
            _843 <= _830;
        4'b1010:
            _843 <= _842;
        default:
            _843 <= _126;
        endcase
    end
    assign _37 = _843;
    always @(posedge _77) begin
        if (_75)
            _126 <= _265;
        else
            _126 <= _37;
    end
    assign _856 = _124 + _806;
    always @* begin
        case (_93)
        4'b1001:
            _858 <= _856;
        default:
            _858 <= _124;
        endcase
    end
    always @* begin
        case (_93)
        4'b1001:
            _853 <= _265;
        default:
            _853 <= _124;
        endcase
    end
    always @* begin
        case (_93)
        4'b1001:
            _849 <= _265;
        default:
            _849 <= _124;
        endcase
    end
    assign _850 = _191 ? _849 : _124;
    assign _854 = _161 ? _853 : _850;
    assign _859 = _131 ? _858 : _854;
    always @* begin
        case (_634)
        4'b1001:
            _845 <= _265;
        default:
            _845 <= _124;
        endcase
    end
    assign _846 = _98 ? _124 : _845;
    assign _847 = _91 ? _124 : _846;
    always @* begin
        case (_85)
        4'b1001:
            _860 <= _847;
        4'b1010:
            _860 <= _859;
        default:
            _860 <= _124;
        endcase
    end
    assign _38 = _860;
    always @(posedge _77) begin
        if (_75)
            _124 <= _265;
        else
            _124 <= _38;
    end
    assign _873 = _122 + _806;
    always @* begin
        case (_93)
        4'b1000:
            _875 <= _873;
        default:
            _875 <= _122;
        endcase
    end
    always @* begin
        case (_93)
        4'b1000:
            _870 <= _265;
        default:
            _870 <= _122;
        endcase
    end
    always @* begin
        case (_93)
        4'b1000:
            _866 <= _265;
        default:
            _866 <= _122;
        endcase
    end
    assign _867 = _191 ? _866 : _122;
    assign _871 = _161 ? _870 : _867;
    assign _876 = _131 ? _875 : _871;
    always @* begin
        case (_634)
        4'b1000:
            _862 <= _265;
        default:
            _862 <= _122;
        endcase
    end
    assign _863 = _98 ? _122 : _862;
    assign _864 = _91 ? _122 : _863;
    always @* begin
        case (_85)
        4'b1001:
            _877 <= _864;
        4'b1010:
            _877 <= _876;
        default:
            _877 <= _122;
        endcase
    end
    assign _39 = _877;
    always @(posedge _77) begin
        if (_75)
            _122 <= _265;
        else
            _122 <= _39;
    end
    assign _890 = _120 + _806;
    always @* begin
        case (_93)
        4'b0111:
            _892 <= _890;
        default:
            _892 <= _120;
        endcase
    end
    always @* begin
        case (_93)
        4'b0111:
            _887 <= _265;
        default:
            _887 <= _120;
        endcase
    end
    always @* begin
        case (_93)
        4'b0111:
            _883 <= _265;
        default:
            _883 <= _120;
        endcase
    end
    assign _884 = _191 ? _883 : _120;
    assign _888 = _161 ? _887 : _884;
    assign _893 = _131 ? _892 : _888;
    always @* begin
        case (_634)
        4'b0111:
            _879 <= _265;
        default:
            _879 <= _120;
        endcase
    end
    assign _880 = _98 ? _120 : _879;
    assign _881 = _91 ? _120 : _880;
    always @* begin
        case (_85)
        4'b1001:
            _894 <= _881;
        4'b1010:
            _894 <= _893;
        default:
            _894 <= _120;
        endcase
    end
    assign _40 = _894;
    always @(posedge _77) begin
        if (_75)
            _120 <= _265;
        else
            _120 <= _40;
    end
    assign _907 = _118 + _806;
    always @* begin
        case (_93)
        4'b0110:
            _909 <= _907;
        default:
            _909 <= _118;
        endcase
    end
    always @* begin
        case (_93)
        4'b0110:
            _904 <= _265;
        default:
            _904 <= _118;
        endcase
    end
    always @* begin
        case (_93)
        4'b0110:
            _900 <= _265;
        default:
            _900 <= _118;
        endcase
    end
    assign _901 = _191 ? _900 : _118;
    assign _905 = _161 ? _904 : _901;
    assign _910 = _131 ? _909 : _905;
    always @* begin
        case (_634)
        4'b0110:
            _896 <= _265;
        default:
            _896 <= _118;
        endcase
    end
    assign _897 = _98 ? _118 : _896;
    assign _898 = _91 ? _118 : _897;
    always @* begin
        case (_85)
        4'b1001:
            _911 <= _898;
        4'b1010:
            _911 <= _910;
        default:
            _911 <= _118;
        endcase
    end
    assign _41 = _911;
    always @(posedge _77) begin
        if (_75)
            _118 <= _265;
        else
            _118 <= _41;
    end
    assign _924 = _116 + _806;
    always @* begin
        case (_93)
        4'b0101:
            _926 <= _924;
        default:
            _926 <= _116;
        endcase
    end
    always @* begin
        case (_93)
        4'b0101:
            _921 <= _265;
        default:
            _921 <= _116;
        endcase
    end
    always @* begin
        case (_93)
        4'b0101:
            _917 <= _265;
        default:
            _917 <= _116;
        endcase
    end
    assign _918 = _191 ? _917 : _116;
    assign _922 = _161 ? _921 : _918;
    assign _927 = _131 ? _926 : _922;
    always @* begin
        case (_634)
        4'b0101:
            _913 <= _265;
        default:
            _913 <= _116;
        endcase
    end
    assign _914 = _98 ? _116 : _913;
    assign _915 = _91 ? _116 : _914;
    always @* begin
        case (_85)
        4'b1001:
            _928 <= _915;
        4'b1010:
            _928 <= _927;
        default:
            _928 <= _116;
        endcase
    end
    assign _42 = _928;
    always @(posedge _77) begin
        if (_75)
            _116 <= _265;
        else
            _116 <= _42;
    end
    assign _941 = _114 + _806;
    always @* begin
        case (_93)
        4'b0100:
            _943 <= _941;
        default:
            _943 <= _114;
        endcase
    end
    always @* begin
        case (_93)
        4'b0100:
            _938 <= _265;
        default:
            _938 <= _114;
        endcase
    end
    always @* begin
        case (_93)
        4'b0100:
            _934 <= _265;
        default:
            _934 <= _114;
        endcase
    end
    assign _935 = _191 ? _934 : _114;
    assign _939 = _161 ? _938 : _935;
    assign _944 = _131 ? _943 : _939;
    always @* begin
        case (_634)
        4'b0100:
            _930 <= _265;
        default:
            _930 <= _114;
        endcase
    end
    assign _931 = _98 ? _114 : _930;
    assign _932 = _91 ? _114 : _931;
    always @* begin
        case (_85)
        4'b1001:
            _945 <= _932;
        4'b1010:
            _945 <= _944;
        default:
            _945 <= _114;
        endcase
    end
    assign _43 = _945;
    always @(posedge _77) begin
        if (_75)
            _114 <= _265;
        else
            _114 <= _43;
    end
    assign _958 = _112 + _806;
    always @* begin
        case (_93)
        4'b0011:
            _960 <= _958;
        default:
            _960 <= _112;
        endcase
    end
    always @* begin
        case (_93)
        4'b0011:
            _955 <= _265;
        default:
            _955 <= _112;
        endcase
    end
    always @* begin
        case (_93)
        4'b0011:
            _951 <= _265;
        default:
            _951 <= _112;
        endcase
    end
    assign _952 = _191 ? _951 : _112;
    assign _956 = _161 ? _955 : _952;
    assign _961 = _131 ? _960 : _956;
    always @* begin
        case (_634)
        4'b0011:
            _947 <= _265;
        default:
            _947 <= _112;
        endcase
    end
    assign _948 = _98 ? _112 : _947;
    assign _949 = _91 ? _112 : _948;
    always @* begin
        case (_85)
        4'b1001:
            _962 <= _949;
        4'b1010:
            _962 <= _961;
        default:
            _962 <= _112;
        endcase
    end
    assign _44 = _962;
    always @(posedge _77) begin
        if (_75)
            _112 <= _265;
        else
            _112 <= _44;
    end
    assign _975 = _110 + _806;
    always @* begin
        case (_93)
        4'b0010:
            _977 <= _975;
        default:
            _977 <= _110;
        endcase
    end
    always @* begin
        case (_93)
        4'b0010:
            _972 <= _265;
        default:
            _972 <= _110;
        endcase
    end
    always @* begin
        case (_93)
        4'b0010:
            _968 <= _265;
        default:
            _968 <= _110;
        endcase
    end
    assign _969 = _191 ? _968 : _110;
    assign _973 = _161 ? _972 : _969;
    assign _978 = _131 ? _977 : _973;
    always @* begin
        case (_634)
        4'b0010:
            _964 <= _265;
        default:
            _964 <= _110;
        endcase
    end
    assign _965 = _98 ? _110 : _964;
    assign _966 = _91 ? _110 : _965;
    always @* begin
        case (_85)
        4'b1001:
            _979 <= _966;
        4'b1010:
            _979 <= _978;
        default:
            _979 <= _110;
        endcase
    end
    assign _45 = _979;
    always @(posedge _77) begin
        if (_75)
            _110 <= _265;
        else
            _110 <= _45;
    end
    assign _992 = _108 + _806;
    always @* begin
        case (_93)
        4'b0001:
            _994 <= _992;
        default:
            _994 <= _108;
        endcase
    end
    always @* begin
        case (_93)
        4'b0001:
            _989 <= _265;
        default:
            _989 <= _108;
        endcase
    end
    always @* begin
        case (_93)
        4'b0001:
            _985 <= _265;
        default:
            _985 <= _108;
        endcase
    end
    assign _986 = _191 ? _985 : _108;
    assign _990 = _161 ? _989 : _986;
    assign _995 = _131 ? _994 : _990;
    always @* begin
        case (_634)
        4'b0001:
            _981 <= _265;
        default:
            _981 <= _108;
        endcase
    end
    assign _982 = _98 ? _108 : _981;
    assign _983 = _91 ? _108 : _982;
    always @* begin
        case (_85)
        4'b1001:
            _996 <= _983;
        4'b1010:
            _996 <= _995;
        default:
            _996 <= _108;
        endcase
    end
    assign _46 = _996;
    always @(posedge _77) begin
        if (_75)
            _108 <= _265;
        else
            _108 <= _46;
    end
    assign _1176 = _106 + _806;
    always @* begin
        case (_93)
        4'b0000:
            _1178 <= _1176;
        default:
            _1178 <= _106;
        endcase
    end
    always @* begin
        case (_93)
        4'b0000:
            _1173 <= _265;
        default:
            _1173 <= _106;
        endcase
    end
    always @* begin
        case (_93)
        4'b0000:
            _1170 <= _265;
        default:
            _1170 <= _106;
        endcase
    end
    assign _1171 = _191 ? _1170 : _106;
    assign _997 = _81 ? _72 : _158;
    always @* begin
        case (_85)
        4'b0001:
            _999 <= _997;
        default:
            _999 <= _158;
        endcase
    end
    assign _47 = _999;
    always @(posedge _77) begin
        if (_75)
            _158 <= _1340;
        else
            _158 <= _47;
    end
    assign _160 = _158 - _640;
    assign _1008 = _155 + _640;
    always @* begin
        case (_93)
        4'b1011:
            _1009 <= _1008;
        default:
            _1009 <= _155;
        endcase
    end
    always @* begin
        case (_93)
        4'b1011:
            _1005 <= _1340;
        default:
            _1005 <= _155;
        endcase
    end
    assign _1006 = _191 ? _1005 : _155;
    assign _1010 = _161 ? _1009 : _1006;
    assign _1011 = _131 ? _155 : _1010;
    always @* begin
        case (_634)
        4'b1011:
            _1001 <= _1340;
        default:
            _1001 <= _155;
        endcase
    end
    assign _1002 = _98 ? _155 : _1001;
    assign _1003 = _91 ? _155 : _1002;
    always @* begin
        case (_85)
        4'b1001:
            _1012 <= _1003;
        4'b1010:
            _1012 <= _1011;
        default:
            _1012 <= _155;
        endcase
    end
    assign _48 = _1012;
    always @(posedge _77) begin
        if (_75)
            _155 <= _1340;
        else
            _155 <= _48;
    end
    assign _1021 = _153 + _640;
    always @* begin
        case (_93)
        4'b1010:
            _1022 <= _1021;
        default:
            _1022 <= _153;
        endcase
    end
    always @* begin
        case (_93)
        4'b1010:
            _1018 <= _1340;
        default:
            _1018 <= _153;
        endcase
    end
    assign _1019 = _191 ? _1018 : _153;
    assign _1023 = _161 ? _1022 : _1019;
    assign _1024 = _131 ? _153 : _1023;
    always @* begin
        case (_634)
        4'b1010:
            _1014 <= _1340;
        default:
            _1014 <= _153;
        endcase
    end
    assign _1015 = _98 ? _153 : _1014;
    assign _1016 = _91 ? _153 : _1015;
    always @* begin
        case (_85)
        4'b1001:
            _1025 <= _1016;
        4'b1010:
            _1025 <= _1024;
        default:
            _1025 <= _153;
        endcase
    end
    assign _49 = _1025;
    always @(posedge _77) begin
        if (_75)
            _153 <= _1340;
        else
            _153 <= _49;
    end
    assign _1034 = _151 + _640;
    always @* begin
        case (_93)
        4'b1001:
            _1035 <= _1034;
        default:
            _1035 <= _151;
        endcase
    end
    always @* begin
        case (_93)
        4'b1001:
            _1031 <= _1340;
        default:
            _1031 <= _151;
        endcase
    end
    assign _1032 = _191 ? _1031 : _151;
    assign _1036 = _161 ? _1035 : _1032;
    assign _1037 = _131 ? _151 : _1036;
    always @* begin
        case (_634)
        4'b1001:
            _1027 <= _1340;
        default:
            _1027 <= _151;
        endcase
    end
    assign _1028 = _98 ? _151 : _1027;
    assign _1029 = _91 ? _151 : _1028;
    always @* begin
        case (_85)
        4'b1001:
            _1038 <= _1029;
        4'b1010:
            _1038 <= _1037;
        default:
            _1038 <= _151;
        endcase
    end
    assign _50 = _1038;
    always @(posedge _77) begin
        if (_75)
            _151 <= _1340;
        else
            _151 <= _50;
    end
    assign _1047 = _149 + _640;
    always @* begin
        case (_93)
        4'b1000:
            _1048 <= _1047;
        default:
            _1048 <= _149;
        endcase
    end
    always @* begin
        case (_93)
        4'b1000:
            _1044 <= _1340;
        default:
            _1044 <= _149;
        endcase
    end
    assign _1045 = _191 ? _1044 : _149;
    assign _1049 = _161 ? _1048 : _1045;
    assign _1050 = _131 ? _149 : _1049;
    always @* begin
        case (_634)
        4'b1000:
            _1040 <= _1340;
        default:
            _1040 <= _149;
        endcase
    end
    assign _1041 = _98 ? _149 : _1040;
    assign _1042 = _91 ? _149 : _1041;
    always @* begin
        case (_85)
        4'b1001:
            _1051 <= _1042;
        4'b1010:
            _1051 <= _1050;
        default:
            _1051 <= _149;
        endcase
    end
    assign _51 = _1051;
    always @(posedge _77) begin
        if (_75)
            _149 <= _1340;
        else
            _149 <= _51;
    end
    assign _1060 = _147 + _640;
    always @* begin
        case (_93)
        4'b0111:
            _1061 <= _1060;
        default:
            _1061 <= _147;
        endcase
    end
    always @* begin
        case (_93)
        4'b0111:
            _1057 <= _1340;
        default:
            _1057 <= _147;
        endcase
    end
    assign _1058 = _191 ? _1057 : _147;
    assign _1062 = _161 ? _1061 : _1058;
    assign _1063 = _131 ? _147 : _1062;
    always @* begin
        case (_634)
        4'b0111:
            _1053 <= _1340;
        default:
            _1053 <= _147;
        endcase
    end
    assign _1054 = _98 ? _147 : _1053;
    assign _1055 = _91 ? _147 : _1054;
    always @* begin
        case (_85)
        4'b1001:
            _1064 <= _1055;
        4'b1010:
            _1064 <= _1063;
        default:
            _1064 <= _147;
        endcase
    end
    assign _52 = _1064;
    always @(posedge _77) begin
        if (_75)
            _147 <= _1340;
        else
            _147 <= _52;
    end
    assign _1073 = _145 + _640;
    always @* begin
        case (_93)
        4'b0110:
            _1074 <= _1073;
        default:
            _1074 <= _145;
        endcase
    end
    always @* begin
        case (_93)
        4'b0110:
            _1070 <= _1340;
        default:
            _1070 <= _145;
        endcase
    end
    assign _1071 = _191 ? _1070 : _145;
    assign _1075 = _161 ? _1074 : _1071;
    assign _1076 = _131 ? _145 : _1075;
    always @* begin
        case (_634)
        4'b0110:
            _1066 <= _1340;
        default:
            _1066 <= _145;
        endcase
    end
    assign _1067 = _98 ? _145 : _1066;
    assign _1068 = _91 ? _145 : _1067;
    always @* begin
        case (_85)
        4'b1001:
            _1077 <= _1068;
        4'b1010:
            _1077 <= _1076;
        default:
            _1077 <= _145;
        endcase
    end
    assign _53 = _1077;
    always @(posedge _77) begin
        if (_75)
            _145 <= _1340;
        else
            _145 <= _53;
    end
    assign _1086 = _143 + _640;
    always @* begin
        case (_93)
        4'b0101:
            _1087 <= _1086;
        default:
            _1087 <= _143;
        endcase
    end
    always @* begin
        case (_93)
        4'b0101:
            _1083 <= _1340;
        default:
            _1083 <= _143;
        endcase
    end
    assign _1084 = _191 ? _1083 : _143;
    assign _1088 = _161 ? _1087 : _1084;
    assign _1089 = _131 ? _143 : _1088;
    always @* begin
        case (_634)
        4'b0101:
            _1079 <= _1340;
        default:
            _1079 <= _143;
        endcase
    end
    assign _1080 = _98 ? _143 : _1079;
    assign _1081 = _91 ? _143 : _1080;
    always @* begin
        case (_85)
        4'b1001:
            _1090 <= _1081;
        4'b1010:
            _1090 <= _1089;
        default:
            _1090 <= _143;
        endcase
    end
    assign _54 = _1090;
    always @(posedge _77) begin
        if (_75)
            _143 <= _1340;
        else
            _143 <= _54;
    end
    assign _1099 = _141 + _640;
    always @* begin
        case (_93)
        4'b0100:
            _1100 <= _1099;
        default:
            _1100 <= _141;
        endcase
    end
    always @* begin
        case (_93)
        4'b0100:
            _1096 <= _1340;
        default:
            _1096 <= _141;
        endcase
    end
    assign _1097 = _191 ? _1096 : _141;
    assign _1101 = _161 ? _1100 : _1097;
    assign _1102 = _131 ? _141 : _1101;
    always @* begin
        case (_634)
        4'b0100:
            _1092 <= _1340;
        default:
            _1092 <= _141;
        endcase
    end
    assign _1093 = _98 ? _141 : _1092;
    assign _1094 = _91 ? _141 : _1093;
    always @* begin
        case (_85)
        4'b1001:
            _1103 <= _1094;
        4'b1010:
            _1103 <= _1102;
        default:
            _1103 <= _141;
        endcase
    end
    assign _55 = _1103;
    always @(posedge _77) begin
        if (_75)
            _141 <= _1340;
        else
            _141 <= _55;
    end
    assign _1112 = _139 + _640;
    always @* begin
        case (_93)
        4'b0011:
            _1113 <= _1112;
        default:
            _1113 <= _139;
        endcase
    end
    always @* begin
        case (_93)
        4'b0011:
            _1109 <= _1340;
        default:
            _1109 <= _139;
        endcase
    end
    assign _1110 = _191 ? _1109 : _139;
    assign _1114 = _161 ? _1113 : _1110;
    assign _1115 = _131 ? _139 : _1114;
    always @* begin
        case (_634)
        4'b0011:
            _1105 <= _1340;
        default:
            _1105 <= _139;
        endcase
    end
    assign _1106 = _98 ? _139 : _1105;
    assign _1107 = _91 ? _139 : _1106;
    always @* begin
        case (_85)
        4'b1001:
            _1116 <= _1107;
        4'b1010:
            _1116 <= _1115;
        default:
            _1116 <= _139;
        endcase
    end
    assign _56 = _1116;
    always @(posedge _77) begin
        if (_75)
            _139 <= _1340;
        else
            _139 <= _56;
    end
    assign _1125 = _137 + _640;
    always @* begin
        case (_93)
        4'b0010:
            _1126 <= _1125;
        default:
            _1126 <= _137;
        endcase
    end
    always @* begin
        case (_93)
        4'b0010:
            _1122 <= _1340;
        default:
            _1122 <= _137;
        endcase
    end
    assign _1123 = _191 ? _1122 : _137;
    assign _1127 = _161 ? _1126 : _1123;
    assign _1128 = _131 ? _137 : _1127;
    always @* begin
        case (_634)
        4'b0010:
            _1118 <= _1340;
        default:
            _1118 <= _137;
        endcase
    end
    assign _1119 = _98 ? _137 : _1118;
    assign _1120 = _91 ? _137 : _1119;
    always @* begin
        case (_85)
        4'b1001:
            _1129 <= _1120;
        4'b1010:
            _1129 <= _1128;
        default:
            _1129 <= _137;
        endcase
    end
    assign _57 = _1129;
    always @(posedge _77) begin
        if (_75)
            _137 <= _1340;
        else
            _137 <= _57;
    end
    assign _1138 = _135 + _640;
    always @* begin
        case (_93)
        4'b0001:
            _1139 <= _1138;
        default:
            _1139 <= _135;
        endcase
    end
    always @* begin
        case (_93)
        4'b0001:
            _1135 <= _1340;
        default:
            _1135 <= _135;
        endcase
    end
    assign _1136 = _191 ? _1135 : _135;
    assign _1140 = _161 ? _1139 : _1136;
    assign _1141 = _131 ? _135 : _1140;
    always @* begin
        case (_634)
        4'b0001:
            _1131 <= _1340;
        default:
            _1131 <= _135;
        endcase
    end
    assign _1132 = _98 ? _135 : _1131;
    assign _1133 = _91 ? _135 : _1132;
    always @* begin
        case (_85)
        4'b1001:
            _1142 <= _1133;
        4'b1010:
            _1142 <= _1141;
        default:
            _1142 <= _135;
        endcase
    end
    assign _58 = _1142;
    always @(posedge _77) begin
        if (_75)
            _135 <= _1340;
        else
            _135 <= _58;
    end
    assign _1158 = _133 + _640;
    always @* begin
        case (_93)
        4'b0000:
            _1160 <= _1158;
        default:
            _1160 <= _133;
        endcase
    end
    always @* begin
        case (_93)
        4'b0000:
            _1155 <= _1340;
        default:
            _1155 <= _133;
        endcase
    end
    assign _1145 = _1144 ? _72 : _188;
    assign _1146 = _81 ? _1145 : _188;
    always @* begin
        case (_85)
        4'b0010:
            _1148 <= _1146;
        default:
            _1148 <= _188;
        endcase
    end
    assign _59 = _1148;
    always @(posedge _77) begin
        if (_75)
            _188 <= _1340;
        else
            _188 <= _59;
    end
    assign _190 = _188 - _640;
    assign _191 = _186 < _190;
    assign _1156 = _191 ? _1155 : _133;
    assign _1161 = _161 ? _1160 : _1156;
    assign _1162 = _131 ? _133 : _1161;
    always @* begin
        case (_634)
        4'b0000:
            _1151 <= _1340;
        default:
            _1151 <= _133;
        endcase
    end
    assign _1152 = _98 ? _133 : _1151;
    assign _1153 = _91 ? _133 : _1152;
    always @* begin
        case (_85)
        4'b0101:
            _1163 <= _1340;
        4'b1001:
            _1163 <= _1153;
        4'b1010:
            _1163 <= _1162;
        default:
            _1163 <= _133;
        endcase
    end
    assign _60 = _1163;
    always @(posedge _77) begin
        if (_75)
            _133 <= _1340;
        else
            _133 <= _60;
    end
    always @* begin
        case (_93)
        0:
            _156 <= _133;
        1:
            _156 <= _135;
        2:
            _156 <= _137;
        3:
            _156 <= _139;
        4:
            _156 <= _141;
        5:
            _156 <= _143;
        6:
            _156 <= _145;
        7:
            _156 <= _147;
        8:
            _156 <= _149;
        9:
            _156 <= _151;
        10:
            _156 <= _153;
        default:
            _156 <= _155;
        endcase
    end
    assign _161 = _156 < _160;
    assign _1174 = _161 ? _1173 : _1171;
    assign _1179 = _131 ? _1178 : _1174;
    assign _634 = _93 + _527;
    always @* begin
        case (_634)
        4'b0000:
            _1166 <= _265;
        default:
            _1166 <= _106;
        endcase
    end
    assign _1167 = _98 ? _106 : _1166;
    assign _1168 = _91 ? _106 : _1167;
    always @* begin
        case (_85)
        4'b0101:
            _1180 <= _265;
        4'b1001:
            _1180 <= _1168;
        4'b1010:
            _1180 <= _1179;
        default:
            _1180 <= _106;
        endcase
    end
    assign _61 = _1180;
    always @(posedge _77) begin
        if (_75)
            _106 <= _265;
        else
            _106 <= _61;
    end
    always @* begin
        case (_93)
        0:
            _129 <= _106;
        1:
            _129 <= _108;
        2:
            _129 <= _110;
        3:
            _129 <= _112;
        4:
            _129 <= _114;
        5:
            _129 <= _116;
        6:
            _129 <= _118;
        7:
            _129 <= _120;
        8:
            _129 <= _122;
        9:
            _129 <= _124;
        10:
            _129 <= _126;
        default:
            _129 <= _128;
        endcase
    end
    assign _131 = _129 < _130;
    assign _1192 = _131 ? _265 : _1190;
    assign _1185 = _89 + _806;
    assign _97 = _95 - _527;
    assign _98 = _93 == _97;
    assign _1183 = _98 ? _89 : _265;
    assign _1186 = _91 ? _1185 : _1183;
    always @* begin
        case (_85)
        4'b0101:
            _1195 <= _265;
        4'b1001:
            _1195 <= _1186;
        4'b1010:
            _1195 <= _1192;
        4'b1101:
            _1195 <= _1194;
        default:
            _1195 <= _89;
        endcase
    end
    assign _62 = _1195;
    always @(posedge _77) begin
        if (_75)
            _89 <= _265;
        else
            _89 <= _62;
    end
    assign _91 = _89 < _90;
    assign _1200 = _91 ? _93 : _1199;
    always @* begin
        case (_85)
        4'b0101:
            _1202 <= _84;
        4'b1001:
            _1202 <= _1200;
        4'b1101:
            _1202 <= _1201;
        default:
            _1202 <= _93;
        endcase
    end
    assign _63 = _1202;
    always @(posedge _77) begin
        if (_75)
            _93 <= _84;
        else
            _93 <= _63;
    end
    always @* begin
        case (_93)
        0:
            _186 <= _163;
        1:
            _186 <= _165;
        2:
            _186 <= _167;
        3:
            _186 <= _169;
        4:
            _186 <= _171;
        5:
            _186 <= _173;
        6:
            _186 <= _175;
        7:
            _186 <= _177;
        8:
            _186 <= _179;
        9:
            _186 <= _181;
        10:
            _186 <= _183;
        default:
            _186 <= _185;
        endcase
    end
    assign _221 = 4'b1101;
    assign _222 = _221 == _85;
    assign _219 = _521 == _85;
    assign _216 = 4'b1011;
    assign _217 = _216 == _85;
    assign _220 = _217 | _219;
    assign _223 = _220 | _222;
    assign _227 = _223 ? _226 : _186;
    assign _238 = _227 + _237;
    assign _1205 = _238[3:0];
    always @* begin
        case (_85)
        4'b0011:
            _1206 <= _1204;
        default:
            _1206 <= _1205;
        endcase
    end
    assign _64 = _1206;
    assign _341 = _340[_64];
    always @(posedge _77) begin
        _342 <= _341;
    end
    assign _1318 = _342 & _626;
    assign _1320 = _1318 == _1349;
    assign _1321 = ~ _1320;
    assign _1352 = _1321 | _1351;
    assign _1355 = _1352 | _1354;
    assign _1356 = _1355 ? _198 : _104;
    assign _87 = 4'b0101;
    assign _1313 = _1301 ? _87 : _85;
    assign _1314 = _264 ? _85 : _1313;
    assign _1312 = _1208 ? _597 : _85;
    assign _1309 = _1280 ? _516 : _85;
    assign _1303 = _245 + _806;
    assign _1300 = 3'b101;
    assign _1301 = _245 == _1300;
    assign _1304 = _1301 ? _245 : _1303;
    assign _1212 = _95 + _527;
    assign _1213 = _264 ? _1212 : _95;
    assign _1210 = _1208 ? _84 : _95;
    always @* begin
        case (_85)
        4'b0011:
            _1214 <= _1210;
        4'b0100:
            _1214 <= _1213;
        default:
            _1214 <= _95;
        endcase
    end
    assign _65 = _1214;
    always @(posedge _77) begin
        if (_75)
            _95 <= _84;
        else
            _95 <= _65;
    end
    assign _263 = _95 < _521;
    assign _1222 = _257 - _640;
    always @* begin
        case (_245)
        3'b101:
            _1224 <= _1222;
        default:
            _1224 <= _257;
        endcase
    end
    assign _1225 = _264 ? _1224 : _257;
    always @* begin
        case (_1216)
        3'b101:
            _1218 <= _72;
        default:
            _1218 <= _257;
        endcase
    end
    assign _1219 = _1144 ? _257 : _1218;
    assign _1220 = _81 ? _1219 : _257;
    always @* begin
        case (_85)
        4'b0010:
            _1226 <= _1220;
        4'b0100:
            _1226 <= _1225;
        default:
            _1226 <= _257;
        endcase
    end
    assign _66 = _1226;
    always @(posedge _77) begin
        if (_75)
            _257 <= _1340;
        else
            _257 <= _66;
    end
    assign _1232 = _255 - _640;
    always @* begin
        case (_245)
        3'b100:
            _1234 <= _1232;
        default:
            _1234 <= _255;
        endcase
    end
    assign _1235 = _264 ? _1234 : _255;
    always @* begin
        case (_1216)
        3'b100:
            _1228 <= _72;
        default:
            _1228 <= _255;
        endcase
    end
    assign _1229 = _1144 ? _255 : _1228;
    assign _1230 = _81 ? _1229 : _255;
    always @* begin
        case (_85)
        4'b0010:
            _1236 <= _1230;
        4'b0100:
            _1236 <= _1235;
        default:
            _1236 <= _255;
        endcase
    end
    assign _67 = _1236;
    always @(posedge _77) begin
        if (_75)
            _255 <= _1340;
        else
            _255 <= _67;
    end
    assign _1242 = _253 - _640;
    always @* begin
        case (_245)
        3'b011:
            _1244 <= _1242;
        default:
            _1244 <= _253;
        endcase
    end
    assign _1245 = _264 ? _1244 : _253;
    always @* begin
        case (_1216)
        3'b011:
            _1238 <= _72;
        default:
            _1238 <= _253;
        endcase
    end
    assign _1239 = _1144 ? _253 : _1238;
    assign _1240 = _81 ? _1239 : _253;
    always @* begin
        case (_85)
        4'b0010:
            _1246 <= _1240;
        4'b0100:
            _1246 <= _1245;
        default:
            _1246 <= _253;
        endcase
    end
    assign _68 = _1246;
    always @(posedge _77) begin
        if (_75)
            _253 <= _1340;
        else
            _253 <= _68;
    end
    assign _1252 = _251 - _640;
    always @* begin
        case (_245)
        3'b010:
            _1254 <= _1252;
        default:
            _1254 <= _251;
        endcase
    end
    assign _1255 = _264 ? _1254 : _251;
    always @* begin
        case (_1216)
        3'b010:
            _1248 <= _72;
        default:
            _1248 <= _251;
        endcase
    end
    assign _1249 = _1144 ? _251 : _1248;
    assign _1250 = _81 ? _1249 : _251;
    always @* begin
        case (_85)
        4'b0010:
            _1256 <= _1250;
        4'b0100:
            _1256 <= _1255;
        default:
            _1256 <= _251;
        endcase
    end
    assign _69 = _1256;
    always @(posedge _77) begin
        if (_75)
            _251 <= _1340;
        else
            _251 <= _69;
    end
    assign _1262 = _249 - _640;
    always @* begin
        case (_245)
        3'b001:
            _1264 <= _1262;
        default:
            _1264 <= _249;
        endcase
    end
    assign _1265 = _264 ? _1264 : _249;
    always @* begin
        case (_1216)
        3'b001:
            _1258 <= _72;
        default:
            _1258 <= _249;
        endcase
    end
    assign _1259 = _1144 ? _249 : _1258;
    assign _1260 = _81 ? _1259 : _249;
    always @* begin
        case (_85)
        4'b0010:
            _1266 <= _1260;
        4'b0100:
            _1266 <= _1265;
        default:
            _1266 <= _249;
        endcase
    end
    assign _70 = _1266;
    always @(posedge _77) begin
        if (_75)
            _249 <= _1340;
        else
            _249 <= _70;
    end
    assign _1272 = _247 - _640;
    always @* begin
        case (_245)
        3'b000:
            _1274 <= _1272;
        default:
            _1274 <= _247;
        endcase
    end
    assign _1275 = _264 ? _1274 : _247;
    assign _72 = s_tdata;
    assign _1215 = 3'b010;
    assign _1216 = _245 - _1215;
    always @* begin
        case (_1216)
        3'b000:
            _1268 <= _72;
        default:
            _1268 <= _247;
        endcase
    end
    assign _1269 = _1144 ? _247 : _1268;
    assign _1270 = _81 ? _1269 : _247;
    always @* begin
        case (_85)
        4'b0010:
            _1276 <= _1270;
        4'b0100:
            _1276 <= _1275;
        default:
            _1276 <= _247;
        endcase
    end
    assign _73 = _1276;
    always @(posedge _77) begin
        if (_75)
            _247 <= _1340;
        else
            _247 <= _73;
    end
    always @* begin
        case (_245)
        0:
            _258 <= _247;
        1:
            _258 <= _249;
        2:
            _258 <= _251;
        3:
            _258 <= _253;
        4:
            _258 <= _255;
        default:
            _258 <= _257;
        endcase
    end
    assign _260 = _258 == _1340;
    assign _261 = ~ _260;
    assign _264 = _261 & _263;
    assign _1305 = _264 ? _245 : _1304;
    assign _1207 = 4'b1111;
    assign _75 = clear;
    assign _77 = clock;
    assign _1286 = _1204 + _527;
    assign _1287 = _1208 ? _1204 : _1286;
    assign _1282 = _1280 ? _84 : _1204;
    assign _1283 = _1278 ? _1204 : _1282;
    assign _1284 = _81 ? _1283 : _1204;
    always @* begin
        case (_85)
        4'b0010:
            _1288 <= _1284;
        4'b0011:
            _1288 <= _1287;
        default:
            _1288 <= _1204;
        endcase
    end
    assign _78 = _1288;
    always @(posedge _77) begin
        if (_75)
            _1204 <= _84;
        else
            _1204 <= _78;
    end
    assign _1208 = _1204 == _1207;
    assign _1299 = _1208 ? _265 : _245;
    assign _1144 = _245 == _806;
    assign _1294 = _1144 ? _1215 : _245;
    assign _1292 = _245 + _806;
    assign _1280 = _245 == _130;
    assign _1295 = _1280 ? _1294 : _1292;
    assign _1296 = _1278 ? _1294 : _1295;
    assign _1297 = _81 ? _1296 : _245;
    assign _1290 = _81 ? _806 : _245;
    always @* begin
        case (_85)
        4'b0001:
            _1306 <= _1290;
        4'b0010:
            _1306 <= _1297;
        4'b0011:
            _1306 <= _1299;
        4'b0100:
            _1306 <= _1305;
        default:
            _1306 <= _245;
        endcase
    end
    assign _79 = _1306;
    always @(posedge _77) begin
        if (_75)
            _245 <= _265;
        else
            _245 <= _79;
    end
    assign _1278 = _245 == _806;
    assign _1310 = _1278 ? _85 : _1309;
    assign _1311 = _81 ? _1310 : _85;
    assign _81 = s_tvalid;
    assign _1308 = _81 ? _604 : _85;
    always @* begin
        case (_85)
        4'b0000:
            _1365 <= _527;
        4'b0001:
            _1365 <= _1308;
        4'b0010:
            _1365 <= _1311;
        4'b0011:
            _1365 <= _1312;
        4'b0100:
            _1365 <= _1314;
        4'b0101:
            _1365 <= _602;
        4'b0110:
            _1365 <= _598;
        4'b0111:
            _1365 <= _436;
        4'b1000:
            _1365 <= _1356;
        4'b1001:
            _1365 <= _1358;
        4'b1010:
            _1365 <= _1362;
        4'b1011:
            _1365 <= _521;
        4'b1100:
            _1365 <= _221;
        4'b1101:
            _1365 <= _1363;
        4'b1110:
            _1365 <= _1364;
        default:
            _1365 <= _85;
        endcase
    end
    assign _82 = _1365;
    always @(posedge _77) begin
        if (_75)
            _85 <= _84;
        else
            _85 <= _82;
    end
    assign _1366 = _527 == _85;
    assign _1368 = _1366 | _1367;
    assign s_tready = _1368;
    assign m_tvalid = _214;
    assign m_tlast = _213;
    assign m_tdata = _211;

endmodule
module range_finder_top (
    m_tready,
    s_tdata,
    s_tvalid,
    clear,
    clock,
    s_tready,
    m_tvalid,
    m_tlast,
    m_tdata
);

    input m_tready;
    input [7:0] s_tdata;
    input s_tvalid;
    input clear;
    input clock;
    output s_tready;
    output m_tvalid;
    output m_tlast;
    output [7:0] m_tdata;

    wire [7:0] _16;
    wire _17;
    wire _18;
    wire _5;
    wire [7:0] _7;
    wire _9;
    wire _11;
    wire _13;
    wire [10:0] _15;
    wire _19;
    assign _16 = _15[10:3];
    assign _17 = _15[2:2];
    assign _18 = _15[1:1];
    assign _5 = m_tready;
    assign _7 = s_tdata;
    assign _9 = s_tvalid;
    assign _11 = clear;
    assign _13 = clock;
    day_12_solver
        day_12_solver
        ( .clock(_13),
          .clear(_11),
          .s_tvalid(_9),
          .s_tdata(_7),
          .m_tready(_5),
          .s_tready(_15[0:0]),
          .m_tvalid(_15[1:1]),
          .m_tlast(_15[2:2]),
          .m_tdata(_15[10:3]) );
    assign _19 = _15[0:0];
    assign s_tready = _19;
    assign m_tvalid = _18;
    assign m_tlast = _17;
    assign m_tdata = _16;

endmodule

// Tiny Tapeout wrapper module
module tt_um_range_finder (
    input  wire       clk,
    input  wire       rst_n,
    input  wire [7:0] ui,
    output wire [7:0] uo,
    inout  wire [7:0] uio
);
    
    // Map Tiny Tapeout pins to day_12_solver interface
    wire clock = clk;
    wire clear = ~rst_n;
    wire s_tvalid = ui[0];
    wire m_tready = ui[1];
    wire [7:0] s_tdata = ui[7:0];
    
    wire s_tready;
    wire m_tvalid;
    wire m_tlast;
    wire [7:0] m_tdata;
    
    // Instantiate the solver
    day_12_solver solver (
        .clock(clock),
        .clear(clear),
        .s_tvalid(s_tvalid),
        .s_tdata(s_tdata),
        .m_tready(m_tready),
        .s_tready(s_tready),
        .m_tvalid(m_tvalid),
        .m_tlast(m_tlast),
        .m_tdata(m_tdata)
    );
    
    // Output mapping
    assign uo[7:0] = m_tdata[7:0];
    
    // Bidirectional mapping
    assign uio[0] = s_tready;
    assign uio[1] = m_tvalid;
    assign uio[2] = m_tlast;
    assign uio[7:3] = 5'b0;

endmodule
